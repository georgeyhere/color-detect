//
//
//
//
`ifndef display_definitions
`define display_definitions
	`define RGB_RED    24'hb71234
	`define RGB_ORNGE  24'hff5800
	`define RGB_YLLW   24'hffd500
	`define RGB_GRN    24'h009b48 
	`define RGB_BLU    24'h0046ad
   
	`define RGB_WHT    24'hffffff
	`define RGB_BLK    24'h0
`endif