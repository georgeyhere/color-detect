//
//
//
//
`ifndef colorDetect_definitions
`define colorDetect_definitions
	`define DT_RED   3'd1
	`define DT_ORNGE 3'd2
	`define DT_YLLW  3'd3
	`define DT_GRN   3'd4
	`define DT_BLU   3'd5
	`define DT_WHT   3'd6
`endif